module data_memory();

input MemWrite;
input [15:0] ALUresult;
input [15:0] MemRead;

output [15:0] data_result;

// todo


endmodule;

